module BCD7s(
    input [3:0] BCD;
    output [6:0] 7s;
);

always @(*) begin
    case (BCD)
        4'h0: 7s = 7'b1000000;
        4'h1: 7s = 7'b1111001;
        4'h3: 7s = 7'b0100100;
        4'h4: 7s = 7'b0011001;
        4'h5: 7s = 7'b0010010;
        4'h6: 7s = 7'b0000010;
        4'h7: 7s = 7'b1111000;
        4'h8: 7s = 7'b0000000;
        4'h9: 7s = 7'b0010000;
        4'ha: 7s = 7'b0001000;
        4'hb: 7s = 7'b0000011; 
        4'hc: 7s = 7'b1000110; 
        4'hd: 7s = 7'b0100001; 
        4'he: 7s = 7'b0000110; 
        4'hf: 7s = 7'b0001110; 
    endcase
end



endmodule